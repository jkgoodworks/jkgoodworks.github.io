--------------------------------------------------------------------------------
--                                  fp32flo
--                    (InputIEEE_8_23_to_8_23_Freq50_uid2)
-- VHDL generated for Zynq7000 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 0.000000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity fp32flo is
    port (clk : in std_logic;
          X : in  std_logic_vector(31 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of fp32flo is
signal expX :  std_logic_vector(7 downto 0);
   -- timing of expX: (c0, 0.000000ns)
signal fracX :  std_logic_vector(22 downto 0);
   -- timing of fracX: (c0, 0.000000ns)
signal sX :  std_logic;
   -- timing of sX: (c0, 0.000000ns)
signal expZero :  std_logic;
   -- timing of expZero: (c0, 0.000000ns)
signal expInfty :  std_logic;
   -- timing of expInfty: (c0, 0.000000ns)
signal fracZero :  std_logic;
   -- timing of fracZero: (c0, 0.000000ns)
signal reprSubNormal :  std_logic;
   -- timing of reprSubNormal: (c0, 0.000000ns)
signal sfracX :  std_logic_vector(22 downto 0);
   -- timing of sfracX: (c0, 0.000000ns)
signal fracR :  std_logic_vector(22 downto 0);
   -- timing of fracR: (c0, 0.000000ns)
signal expR :  std_logic_vector(7 downto 0);
   -- timing of expR: (c0, 0.000000ns)
signal infinity :  std_logic;
   -- timing of infinity: (c0, 0.000000ns)
signal zero :  std_logic;
   -- timing of zero: (c0, 0.000000ns)
signal NaN :  std_logic;
   -- timing of NaN: (c0, 0.000000ns)
signal exnR :  std_logic_vector(1 downto 0);
   -- timing of exnR: (c0, 0.000000ns)
begin
   expX  <= X(30 downto 23);
   fracX  <= X(22 downto 0);
   sX  <= X(31);
   expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
   expInfty  <= '1' when expX = (7 downto 0 => '1') else '0';
   fracZero <= '1' when fracX = (22 downto 0 => '0') else '0';
   reprSubNormal <= fracX(22);
   -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
   -- we can represent subnormal numbers whose mantissa field begins with a 1
   sfracX <= fracX(21 downto 0) & '0' when (expZero='1' and reprSubNormal='1')    else fracX;
   fracR <= sfracX;
   -- copy exponent. This will be OK even for subnormals, zero and infty since in such cases the exn bits will prevail
   expR <= expX;
   infinity <= expInfty and fracZero;
   zero <= expZero and not reprSubNormal;
   NaN <= expInfty and not fracZero;
   exnR <= 
           "00" when zero='1' 
      else "10" when infinity='1' 
      else "11" when NaN='1' 
      else "01" ;  -- normal number
   R <= exnR & sX & expR & fracR; 
end architecture;

